parameter DATA_WORDS = 0;
