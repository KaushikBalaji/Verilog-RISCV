parameter INSTR_WORDS = 21;
