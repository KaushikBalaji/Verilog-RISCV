parameter DATA_WORDS = 1;
