`ifndef INSTR_SIZE_VH
`define INSTR_SIZE_VH

`define INSTR_WORDS 6

`endif
