parameter INSTR_WORDS = 5;
